/* ECPE 174 - Adv. Digital Design 
	Lab #  : 
	Author : Kelvin Flores 
	Date : 
	Due :  
	
*/

module vgaSync(		input logic clock,
							input logic button,
							output logic );


	
endmodule
						  
						  