library verilog;
use verilog.vl_types.all;
entity testGrid is
end testGrid;
