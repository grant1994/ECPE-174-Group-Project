library verilog;
use verilog.vl_types.all;
entity TB_mem512 is
end TB_mem512;
