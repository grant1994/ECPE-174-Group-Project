library verilog;
use verilog.vl_types.all;
entity TB_mem64 is
end TB_mem64;
