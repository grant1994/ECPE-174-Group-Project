/* ECPE 174 - Adv. Digital Design 
	Lab #  : 
	Author : Kelvin Flores 
	Date : 
	Due :  
	
*/

module XXXXXX (input logic clock,
						  input logic ,
						  output logic );


	
endmodule
						  
						  