/* ECPE 174 - Adv. Digital Design 
	Lab #  : 
	Author : Kelvin Flores 
	Date : 
	Due :  
	
*/

`timescale 1ns/1ns
module ####();
  
	logic clock = 1'b0;

	always #25 clock <= ~clock;
	
	
	
  initial
  begin

     
  end

  
endmodule