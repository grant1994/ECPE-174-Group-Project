library verilog;
use verilog.vl_types.all;
entity testCompare is
end testCompare;
