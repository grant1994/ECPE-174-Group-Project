library verilog;
use verilog.vl_types.all;
entity TB_playGame is
end TB_playGame;
