library verilog;
use verilog.vl_types.all;
entity TB_draw is
end TB_draw;
