library verilog;
use verilog.vl_types.all;
entity TB_arrowKeys is
end TB_arrowKeys;
