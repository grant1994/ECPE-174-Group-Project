library verilog;
use verilog.vl_types.all;
entity TB_dpm is
end TB_dpm;
